`timescale 1ns/1ps
`define MEM_DEPTH  1024
`define MEM_WIDTH  8
`define WORD_WIDTH 16
`define CLOCK_PD 20

`include "winnerPolicy.v"

module tb_winnerPolicy();
    reg clock, nreset;
endmodule