module winnerPolicy(clock, reset, v)